* Brown-out Threshold Analysis
* ============================
* Determines the minimum AC input voltage where MCU supply stays stable
* Uses slow ramp-down to find threshold without transient effects
*
* Key questions:
*   1. At what AC RMS voltage does 12V rail enter dropout?
*   2. At what AC RMS voltage does 3.3V rail fall below BOR?
*   3. What safety margin exists at nominal 120V?

.title Softstart MCU Supply - Brown-out Threshold Analysis

* Include component models
.include lib/components.lib

*=============================================================================
* Circuit Parameters
*=============================================================================

.param GEN_FREQ=60
.param GEN_ZINT=2

* Voltage ramp parameters
.param V_START=120           ; Start at nominal
.param V_END=40              ; Ramp down to find threshold
.param RAMP_TIME=5           ; Slow ramp to avoid transients

* MCU load current (worst case)
.param MCU_ILOAD=50m         ; 50mA worst case

*=============================================================================
* Power Source - Ramping Generator
*=============================================================================

* Ramp control (120V RMS down to 40V RMS over RAMP_TIME)
Vctrl ramp_ctrl 0 PWL(0 {V_START} {RAMP_TIME} {V_END})

* Peak voltage tracks RMS
Bgen ac_hot_int 0 V={sin(6.28318 * GEN_FREQ * time) * V(ramp_ctrl) * 1.414}
Rgen ac_hot_int ac_l {GEN_ZINT}

Vn ac_n 0 0

*=============================================================================
* MCU Power Supply Chain
*=============================================================================

* Bridge rectifier
D1 ac_l rect_pos DFAST
D2 ac_n rect_pos DFAST
D3 0 ac_l DFAST
D4 0 ac_n DFAST
.model DFAST D(Is=1e-14 Rs=0.1 BV=600)

* Bulk capacitor C8 (1000uF)
C_bulk rect_pos 0 1000u IC=170

* LM7812
Xlm7812 rect_pos 0 rail_12v LM7812

* C9 (10uF)
C9 rail_12v 0 10u IC=12

* AMS1117-3.3
Xams1117 rail_12v 0 rail_3v3 AMS1117

* Output caps
C1 rail_3v3 0 10u IC=3.3
C2 rail_3v3 0 10u IC=3.3

* MCU load (worst case current draw)
Rmcu rail_3v3 0 {3.3/MCU_ILOAD}

*=============================================================================
* Additional Loads on 12V Rail
*=============================================================================

* Gate drivers (4x UCC27511A, ~1mA each quiescent, up to 10mA switching)
Rgate_drivers rail_12v 0 {12/0.04}

* Status LED (~10mA)
Rled rail_12v 0 {12/0.01}

*=============================================================================
* Threshold Detection
*=============================================================================

* 12V dropout indicator (1 when rail < 11V)
B12v_dropout 12v_dropout 0 V={3.3 * (V(rail_12v) < 11 ? 1 : 0)}

* 3.3V BOR indicator (1 when rail < 2.0V)
B3v3_bor 3v3_bor 0 V={3.3 * (V(rail_3v3) < 2.0 ? 1 : 0)}

* 3.3V warning indicator (1 when rail < 3.0V)
B3v3_warn 3v3_warn 0 V={3.3 * (V(rail_3v3) < 3.0 ? 1 : 0)}

*=============================================================================
* Analysis
*=============================================================================

.tran 1m {RAMP_TIME} 0 1m

*=============================================================================
* Output Control
*=============================================================================

.control
    run

    set hcopydevtype=svg

    * Plot 1: Input vs output voltages
    plot v(ramp_ctrl) v(rect_pos)/2 v(rail_12v) v(rail_3v3)*5 title 'Supply Rails vs AC Input'
    + xlabel 'Time (s)' ylabel 'Voltage (V)'

    * Plot 2: Threshold indicators
    plot v(ramp_ctrl) v(12v_dropout)*30 v(3v3_warn)*30 v(3v3_bor)*30 title 'Threshold Crossings'
    + xlabel 'Time (s)' ylabel 'V_RMS / Indicator'

    * Plot 3: Zoom on regulation limits
    plot v(rail_12v) v(rail_3v3)*3 title '12V and 3.3V Rails (3.3V scaled 3x)'
    + xlabel 'Time (s)' ylabel 'Voltage (V)'

    * Measurements - find when each threshold is crossed
    echo ""
    echo "=== Brown-out Threshold Measurements ==="

    * Find AC voltage when 12V drops below 11V (regulation limit)
    meas tran t_12v_dropout WHEN v(rail_12v)=11 FALL=1
    if t_12v_dropout > 0
        meas tran vac_12v_dropout FIND v(ramp_ctrl) AT=t_12v_dropout
        echo "12V rail dropout (< 11V) at AC RMS: $&vac_12v_dropout V"
    end

    * Find AC voltage when 3.3V drops below 3.0V (warning)
    meas tran t_3v3_warn WHEN v(rail_3v3)=3.0 FALL=1
    if t_3v3_warn > 0
        meas tran vac_3v3_warn FIND v(ramp_ctrl) AT=t_3v3_warn
        echo "3.3V rail warning (< 3.0V) at AC RMS: $&vac_3v3_warn V"
    end

    * Find AC voltage when 3.3V drops below 2.0V (BOR)
    meas tran t_3v3_bor WHEN v(rail_3v3)=2.0 FALL=1
    if t_3v3_bor > 0
        meas tran vac_3v3_bor FIND v(ramp_ctrl) AT=t_3v3_bor
        echo "3.3V rail BOR (< 2.0V) at AC RMS: $&vac_3v3_bor V"
    end

    * Calculate margins
    echo ""
    echo "=== Safety Margins at 120V RMS ==="

    meas tran v12v_at_120 FIND v(rail_12v) AT=0.1
    meas tran v3v3_at_120 FIND v(rail_3v3) AT=0.1
    echo "At 120V AC: 12V rail = $&v12v_at_120 V, 3.3V rail = $&v3v3_at_120 V"

    meas tran v12v_at_90 FIND v(rail_12v) WHEN v(ramp_ctrl)=90
    meas tran v3v3_at_90 FIND v(rail_3v3) WHEN v(ramp_ctrl)=90
    echo "At 90V AC (25% droop): 12V rail = $&v12v_at_90 V, 3.3V rail = $&v3v3_at_90 V"

    * Minimum AC voltage for stable operation
    echo ""
    echo "=== Minimum Operating Voltage ==="
    if t_3v3_bor > 0
        echo "MCU brown-out occurs at AC RMS: $&vac_3v3_bor V"
        let margin = 120 - vac_3v3_bor
        echo "Safety margin from 120V nominal: $&margin V RMS"
        let pct_margin = 100 * (120 - vac_3v3_bor) / 120
        echo "Percentage margin: $&pct_margin %"
    else
        echo "MCU stays powered across entire test range (40-120V RMS)"
    end

    * Write data
    wrdata results/brownout_threshold.csv v(ramp_ctrl) v(rect_pos) v(rail_12v) v(rail_3v3)

.endc

.end
